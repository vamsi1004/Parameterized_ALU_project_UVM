`include "defines.svh"
class alu_sequence1 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence1)
  
  function new(string name  = "alu_sequence");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 0;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence2 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence2)
  
  function new(string name  = "alu_sequence2");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 1;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence3 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence3)
  
  function new(string name  = "alu_sequence3");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 2;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence4 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence4)
  
  function new(string name  = "alu_sequence4");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 3;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence5 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence5)
  
  function new(string name  = "alu_sequence5");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 4;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence6 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence6)
  
  function new(string name  = "alu_sequence6");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 5;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence7 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence7)
  
  function new(string name  = "alu_sequence7");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 6;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence8 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence8)
  
  function new(string name  = "alu_sequence8");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 7;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence9 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence9)
  
  function new(string name  = "alu_sequence9");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 8;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence10 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence10)
  
  function new(string name  = "alu_sequence10");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD ==9;MODE == 1;INP_VALID == 3;})
  endtask 
endclass 

class alu_sequence11 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence11)
  
  function new(string name  = "alu_sequence10");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD ==10;MODE == 1;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence12 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence12)
  
  function new(string name  = "alu_sequence10");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD ==0;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence13 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence13)
  
  function new(string name  = "alu_sequence13");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD ==1;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence14 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence14)
  
  function new(string name  = "alu_sequence14");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 2;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence15 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence15)
  
  function new(string name  = "alu_sequence15");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 3;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence16 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence16)
  
  function new(string name  = "alu_sequence16");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 4;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence17 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence17)
  
  function new(string name  = "alu_sequence17");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 5;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence18 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence18)
  
  function new(string name  = "alu_sequence18");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 6;MODE == 0;})
  endtask 
endclass

class alu_sequence19 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence19)
  
  function new(string name  = "alu_sequence19");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 7;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence20 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence20)
  
  function new(string name  = "alu_sequence20");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 8;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence21 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence21)
  
  function new(string name  = "alu_sequence21");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 9;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence22 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence22)
  
  function new(string name  = "alu_sequence22");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 10;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence23 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence23)
  
  function new(string name  = "alu_sequence23");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 11;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence24 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence24)
  
  function new(string name  = "alu_sequence24");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 12;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence25 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence25)
  
  function new(string name  = "alu_sequence25");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 13;MODE == 0;INP_VALID == 3;})
  endtask 
endclass

class alu_sequence26 extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(alu_sequence26)
  
  function new(string name  = "alu_sequence26");
    super.new(name);
  endfunction 
  
  virtual task body();
    req = alu_seq_item::type_id::create("req");
    `uvm_rand_send_with(req,{CMD == 0;MODE == 1;INP_VALID == 2;})
  endtask 
endclass


class virtual_sequence extends uvm_sequence #(alu_seq_item);
  
  `uvm_object_utils(virtual_sequence)
  
  alu_sequence1 seq1;
  alu_sequence2 seq2;
  alu_sequence3 seq3;
  alu_sequence4 seq4;
  alu_sequence5 seq5;
  alu_sequence6 seq6;
  alu_sequence7 seq7;
  alu_sequence8 seq8;
  alu_sequence9 seq9;
  alu_sequence10 seq10;
  alu_sequence11 seq11;
  alu_sequence12 seq12;
  alu_sequence13 seq13;
  alu_sequence14 seq14;
  alu_sequence15 seq15;
  alu_sequence16 seq16;
  alu_sequence17 seq17;
  alu_sequence18 seq18;
  alu_sequence19 seq19;
  alu_sequence20 seq20;
  alu_sequence21 seq21;
  alu_sequence22 seq22;
  alu_sequence23 seq23;
  alu_sequence24 seq24;
  alu_sequence25 seq25;
  alu_sequence26 seq26;
  
  alu_sequencer seqA;
  
  function new(string name = "v_seq");
    super.new(name);
  endfunction 
  
  virtual task body();
    seq1 = alu_sequence1::type_id::create("seq1");
    seq2 = alu_sequence2::type_id::create("seq2");
    seq3 = alu_sequence3::type_id::create("seq3");
    seq4 = alu_sequence4::type_id::create("seq4");
    seq5 = alu_sequence5::type_id::create("seq5");
    seq6 = alu_sequence6::type_id::create("seq6");
    seq7 = alu_sequence7::type_id::create("seq7");
    seq8 = alu_sequence8::type_id::create("seq8");
    seq9 = alu_sequence9::type_id::create("seq9");
    seq10 = alu_sequence10::type_id::create("seq10");
    seq11 = alu_sequence11::type_id::create("seq11");
    seq12 = alu_sequence12::type_id::create("seq12");
    seq13 = alu_sequence13::type_id::create("seq13");
    seq14 = alu_sequence14::type_id::create("seq14");
    seq15 = alu_sequence15::type_id::create("seq15");
    seq16 = alu_sequence16::type_id::create("seq16");
    seq17 = alu_sequence17::type_id::create("seq17");
    seq18 = alu_sequence18::type_id::create("seq18");
    seq19 = alu_sequence19::type_id::create("seq19");
    seq20 = alu_sequence20::type_id::create("seq20");
    seq21 = alu_sequence21::type_id::create("seq21");
    seq22 = alu_sequence22::type_id::create("seq22");
    seq23 = alu_sequence23::type_id::create("seq23");
    seq24 = alu_sequence24::type_id::create("seq24");
    seq25 = alu_sequence25::type_id::create("seq25");
    seq26 = alu_sequence26::type_id::create("seq26");
    
    seq1.start(seqA);
    seq2.start(seqA);
    seq3.start(seqA);
    seq4.start(seqA);
    seq5.start(seqA);
    seq6.start(seqA);
    seq7.start(seqA);
    seq8.start(seqA);
    seq9.start(seqA);
    seq10.start(seqA);
    seq11.start(seqA);
    seq12.start(seqA);
    seq13.start(seqA);
    seq14.start(seqA);
    seq15.start(seqA);
    seq16.start(seqA);
    seq17.start(seqA);
    seq18.start(seqA);
    seq19.start(seqA);
    seq20.start(seqA);
    seq21.start(seqA);
    seq22.start(seqA);
    seq23.start(seqA);
    seq24.start(seqA);
    seq25.start(seqA);
    seq26.start(seqA);
  endtask 

endclass

